SIGNAL I_BUFFERED : std_logic_vector(0 TO %%I_MAX);
SIGNAL C_SIG : std_logic_vector(0 TO %%C_MAX);
SIGNAL STATE, NEXTSTATE : std_logic_vector(%%STATEWIDTH_M1 DOWNTO 0);